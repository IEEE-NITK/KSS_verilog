module or_imp(input in_1, //first input to or gate
			   input in_2, //second input to or gate
			   input out); // output of or gate
			   
	assign out = in_1 | in_2;

endmodule	